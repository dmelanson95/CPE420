LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_SIGNED;


ENTITY MIPS_ALU_tb IS
END MIPS_ALU_tb;

ARCHITECTURE Behavior OF MIPS_ALU_tb IS

COMPONENT MIPS_ALU IS
PORT
(

	ALU_CTL : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	A, B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	ALU_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	ZERO : OUT STD_LOGIC
);
END COMPONENT;

SIGNAL ALU_CTL : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL A, B : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL ALU_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL ZERO : STD_LOGIC;

SIGNAL A_VAL : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');			-- DECIMAL 64 --
SIGNAL B_VAL : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');				-- DECIMAL 128 --

BEGIN
	
	UUT: MIPS_ALU PORT MAP (
		ALU_CTL => ALU_CTL,
		A => A,
		B => B,
		ALU_OUT => ALU_OUT,
		ZERO => ZERO
	);
	
	PROCESS
	BEGIN
			-- AND --
			A <= A_VAL;
			B <= B_VAL;
			ALU_CTL <= "0000";
			WAIT FOR 100 NS;
			
			
			-- OR --
			A <= A_VAL;
			B <= B_VAL;
			ALU_CTL <= "0001";
			WAIT FOR 100 NS;
			
			-- ADDITION --
			-- RESULT SHOULD BE SAME AS OR
			A <= A_VAL;
			B <= B_VAL;
			ALU_CTL <="0010";
			WAIT FOR 100 NS;
			
			-- SUBTRACT --
			A <= A_VAL;
			B <= B_VAL;
			ALU_CTL <= "0110";
			WAIT FOR 100 NS;
			
			-- SET ON LESS THAN --
			-- RESULT SHOULD BE 1'S
			A <= A_VAL;
			B <= B_VAL;
			ALU_CTL <="0111";
			WAIT FOR 100 NS;
			
			-- NOR --
			A <= A_VAL;
			B <= B_VAL;
			ALU_CTL <= "1100";
			WAIT FOR 100 NS;
			
	END PROCESS;
	
END Behavior;
