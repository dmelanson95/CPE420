LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_SIGNED;


ENTITY MIPS_ALU IS
PORT
(

	ALU_CTL : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	A, B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	ALU_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	ZERO : OUT STD_LOGIC
);
END MIPS_ALU;

ARCHITECTURE Behavior OF MIPS_ALU IS

SIGNAL ALU_OUT_BUFF : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
	
	PROCESS(ALU_CTL)
		BEGIN
		CASE ALU_CTL IS
			WHEN "0000" =>
				ALU_OUT_BUFF <= A AND B;
				
			WHEN "0001" =>
				ALU_OUT_BUFF <= A OR B;
				
			WHEN "0010" =>
				ALU_OUT_BUFF <= STD_LOGIC_VECTOR(TO_SIGNED((TO_INTEGER(SIGNED(A)) + TO_INTEGER(SIGNED(B))), 32));
				
			WHEN "0110" =>
				ALU_OUT_BUFF <= STD_LOGIC_VECTOR(TO_SIGNED((TO_INTEGER(SIGNED(A)) - TO_INTEGER(SIGNED(B))), 32));
				
			WHEN "0111" =>
				IF A <= B THEN 
					ALU_OUT_BUFF <= (OTHERS => '1');
				ELSE
					ALU_OUT_BUFF <= (OTHERS => '0');
				END IF;
				
			WHEN "1100" =>
				ALU_OUT_BUFF <= A NOR B;
			
			WHEN OTHERS =>
				ALU_OUT_BUFF <= (OTHERS => '0');
				
		END CASE;
	END PROCESS;
	
	PROCESS(ALU_OUT_BUFF) IS
	BEGIN
		IF ALU_OUT_BUFF = "00000000000000000000000000000000" THEN
			ZERO <= '1';
		ELSE
			ZERO <= '0';
		END IF;
	END PROCESS;
	
	ALU_OUT <= ALU_OUT_BUFF;
	
END Behavior;